-------------------------------------------------------------------------------
-- Title      : Interfacing cicuit code
-- Project    : 
-------------------------------------------------------------------------------
-- File       : interface.vhd
-- Author     : Aniket <anktdshmkh@gmail.com>
-- Company    : 
-- Last update: 2006/06/17
-- Platform   : 
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2006/06/14  1.0      V1	Created
-------------------------------------------------------------------------------

entity interface_unit is
  
end interface_unit;

architecture interface_unit_A of interface_unit is

begin  -- interface_unit_A

  

end interface_unit_A;
